library verilog;
use verilog.vl_types.all;
entity ascii_decoder_hex_vlg_vec_tst is
end ascii_decoder_hex_vlg_vec_tst;
